* Mary Had a Little Lamb FSM Subcircuit Definition
.SUBCKT MaryLambFSM_new CLK RST START NOTE2 NOTE1 NOTE0 STATE2 STATE1 STATE0 DONE
* Parameters
.param VDD=5

* State Storage using existing Register components
* Each Register has CLK and D[3:0] inputs, Q[3:0] and Qb[3:0] outputs
* We'll use only one bit from each register for our state bits
X1 CLK D0 Q0 Qb0 dff
X2 CLK D1 Q1 Qb1 dff
X3 CLK D2 Q2 Qb2 dff

* Next State Logic using behavioral sources
* State sequence: 000->001->010->011->100->101->110->111
B_D0 D0 0 V= if(V(RST)>2.5, 0,
               if(V(START)>2.5 & V(Q2,Q1,Q0)==b'000, 1,
               if(V(Q2,Q1,Q0)==b'001, 0,
               if(V(Q2,Q1,Q0)==b'010, 1,
               if(V(Q2,Q1,Q0)==b'011, 0,
               if(V(Q2,Q1,Q0)==b'100, 1,
               if(V(Q2,Q1,Q0)==b'101, 0,
               if(V(Q2,Q1,Q0)==b'110, 1, 0))))))))

B_D1 D1 0 V= if(V(RST)>2.5, 0,
               if(V(START)>2.5 & V(Q2,Q1,Q0)==b'000, 0,
               if(V(Q2,Q1,Q0)==b'001, 1,
               if(V(Q2,Q1,Q0)==b'010, 1,
               if(V(Q2,Q1,Q0)==b'011, 0,
               if(V(Q2,Q1,Q0)==b'100, 0,
               if(V(Q2,Q1,Q0)==b'101, 1,
               if(V(Q2,Q1,Q0)==b'110, 1, 1))))))))

B_D2 D2 0 V= if(V(RST)>2.5, 0,
               if(V(START)>2.5 & V(Q2,Q1,Q0)==b'000, 0,
               if(V(Q2,Q1,Q0)==b'001, 0,
               if(V(Q2,Q1,Q0)==b'010, 0,
               if(V(Q2,Q1,Q0)==b'011, 1,
               if(V(Q2,Q1,Q0)==b'100, 1,
               if(V(Q2,Q1,Q0)==b'101, 1,
               if(V(Q2,Q1,Q0)==b'110, 1, 1))))))))

* Note Output Logic (3=E, 2=D, 1=C, 0=Rest)
B_NOTE2 NOTE2 0 V= if(V(Q2,Q1,Q0)==b'001 | V(Q2,Q1,Q0)==b'101 | V(Q2,Q1,Q0)==b'110, 1, 0)
B_NOTE1 NOTE1 0 V= if(V(Q2,Q1,Q0)==b'010 | V(Q2,Q1,Q0)==b'100, 1, 0)
B_NOTE0 NOTE0 0 V= if(V(Q2,Q1,Q0)==b'011, 1, 0)

* State Output
B_STATE2 STATE2 0 V=V(Q2)
B_STATE1 STATE1 0 V=V(Q1)
B_STATE0 STATE0 0 V=V(Q0)

* Done Signal (active when in state 111)
B_DONE DONE 0 V= if(V(Q2,Q1,Q0)==b'111, {VDD}, 0)

* Pull-down resistors for stability
R1 Q0 0 1k
R2 Q1 0 1k
R3 Q2 0 1k
R4 D0 0 1k
R5 D1 0 1k
R6 D2 0 1k

.ENDS MaryLambFSM_new
